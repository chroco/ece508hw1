
// fulladd4.v - 4-bit binary adder
//
// <your name>
// <date>
//
// Description:
// ------------
// <your description of what the module does>
//
module fulladd4 (
	input logic	[3:0]		a, b,
	input logic				c_in,
	output logic	[3:0]	s,
	output logic			c_out
);

// ADD YOUR CODE HERE

endmodule: fulladd4


