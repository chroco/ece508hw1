


// bcd_adder.v - 4-bit BCD Adder with illegal input detection using Verilog dataflow modeling
//
// <your name>
// <date>
//
// Description:
// ------------
// <your description of what the module does>
//
module bcd_adder (
	input logic	[3:0]		X, Y,
	input logic				c_in,
	output logic			c_out,
	output logic	[7:0]	result,
	output logic			out_of_range
);

// ADD YOUR CODE HERE

endmodule: bcd_adder
